--branch equal control---------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;
entity branch is
  port(rst :in std_logic;
    beq :in std_logic;
    opcode :in std_logic_vector(2 downto 0);
    pccontrol :in std_logic;
    pcen:out std_logic);
  end branch;
  
architecture bhv of branch is 
begin
  process(rst,beq,opcode,pccontrol)
  variable isbeq : std_logic;
  variable gate: std_logic :='0';
  begin
    if(rst = '1') then
       pcen <= '0';
     else
  case opcode is
  when "100" => isbeq:='1';
  when others => isbeq:='0';
  end case;
  if isbeq='1' and beq = '1' then
      gate:='1';
    else
      gate:='0';
  end if;
  pcen<= (gate or pccontrol);
end if;
end process;
end architecture bhv;

--4 to 1 mux-------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity mux4 is
port(rst:in std_logic;
c : in std_logic_vector(31 downto 0);
d : in std_logic_vector(31 downto 0);
e : in std_logic_vector(31 downto 0);
f : in std_logic_vector(31 downto 0);
s : in std_logic_vector(1 downto 0);
muxoutput : out std_logic_vector(31 downto 0));
end mux4;

architecture bhv of mux4 is
begin
process(rst,s,c,d,e,f)
begin
  if(rst = '1') then
  muxoutput <= "00000000000000000000000000000000";
else
case s is
when "00"=> muxoutput <= c;
when "01"=> muxoutput <= d;
when "10"=> muxoutput <= e;
when "11"=> muxoutput <= f;
when others => null;
end case;
end if;
end process;
end bhv;

--random module-------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
entity ram_module is
port(rst :in std_logic;
clk : in std_logic;
enable : in std_logic;
R_W : in std_logic;
addr : in std_logic_vector (31 downto 0);
data_in : in std_logic_vector (31 downto 0);
data_out : out std_logic_vector (31 downto 0));
end ram_module;
--please replace the ram_module with the ram_test file I provided
architecture bhv of ram_module is
type memory is array (0 to 65536) of std_logic_vector(31 downto 0);
signal mem: memory;
begin
process(rst,clk,R_W,addr,enable)
  begin
    if (rst ='1') then
mem(0) <= conv_std_logic_vector(8454155,32);
mem(1) <= conv_std_logic_vector(8519692,32);
mem(2) <= conv_std_logic_vector(8585227,32);
mem(3) <= conv_std_logic_vector(8650765,32);
mem(4) <= conv_std_logic_vector(8716299,32);
mem(5) <= conv_std_logic_vector(17432580,32);
mem(6) <= conv_std_logic_vector(786433,32);
mem(7) <= conv_std_logic_vector(1835011,32);
mem(8) <= conv_std_logic_vector(22347776,32);
mem(9) <= conv_std_logic_vector(29360128,32);
mem(10) <= conv_std_logic_vector(25165824,32);
mem(11) <= conv_std_logic_vector(0,32);
mem(12) <= conv_std_logic_vector(5,32);
mem(13) <= conv_std_logic_vector(1,32); 
data_out <=conv_std_logic_vector(0,32);
else
if(clk'event and clk='1') then
if(enable='1') then
if(R_W='0') then
data_out<=mem(conv_integer(addr));
else
mem(conv_integer(addr))<=data_in;
end if;
end if;
end if;
end if;
end process;
end bhv;

--2 to 1 mux-------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity mux2 is
port(rst: in std_logic;
c : in std_logic_vector(31 downto 0);
d : in std_logic_vector(31 downto 0);
s : in std_logic;
muxoutput : out std_logic_vector(31 downto 0));
end mux2;

architecture bhv of mux2 is
begin
process(rst,s,c,d)
begin
  if(rst ='1') then 
  muxoutput <= "00000000000000000000000000000000";
else
case s is
when '0'=> muxoutput <= c;
when '1'=> muxoutput <= d;
when others => null;
end case;
end if;
end process;
end bhv;

--register mux-----------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity muxr is
port(rst : in std_logic;
c : in std_logic_vector(2 downto 0);
d : in std_logic_vector(2 downto 0);
s : in std_logic;
muxoutput : out std_logic_vector(2 downto 0));
end muxr;

architecture bhv of muxr is
begin
process(rst,s,c,d)
begin
  if(rst ='1') then 
  muxoutput <= "000";
else
case s is
when '0'=> muxoutput <= c;
when '1'=> muxoutput <= d;
when others => null;
end case;
end if;
end process;
end bhv;

--sign extension unit----------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity sext is
port(rst :in std_logic;
A : in std_logic_vector (15 downto 0);
O : out std_logic_vector (31 downto 0));
end sext;

architecture bhv of sext is
begin
process(A,rst)
begin
  if(rst = '1') then
     O<= "00000000000000000000000000000000";
   else
if (A(15) = '1') then
O <= "1111111111111111" & A;
elsif (A(15) = '0') then
O <= "0000000000000000" & A;
end if;
end if;
end process;
end bhv;

--32 bit register--------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
entity reg is
  port(rst: in std_logic;
clk : in std_logic;
enable : in std_logic;
data : in std_logic_vector (31 downto 0);
O : out std_logic_vector (31 downto 0));
end reg;

architecture bhv of reg is
begin
process(rst,clk,enable)
variable temp:std_logic_vector (31 downto 0):="00000000000000000000000000000000";
begin
  if (rst ='1') then
    O<="00000000000000000000000000000000";
  else
if (clk'event and clk='1') then
if enable='1' then
O<=data;
temp:=data;
else
O<=temp;
end if;
end if;
end if;
end process;
end bhv;

--8x32 register bank-----------------------------
LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
entity register_file is
port(rst : in std_logic;
clk : in std_logic;
DR_enable : in std_logic;
DR_address : in std_logic_vector (2 downto 0);
SR1_address: in std_logic_vector(2 downto 0);
SR2_address: in std_logic_vector(2 downto 0);
data_in: in std_logic_vector (31 downto 0);
SR1_out: out std_logic_vector (31 downto 0);
SR2_out: out std_logic_vector (31 downto 0);
r0: out std_logic_vector(31 downto 0);
r1: out std_logic_vector(31 downto 0);
r2: out std_logic_vector(31 downto 0);
r3: out std_logic_vector(31 downto 0);
r4: out std_logic_vector(31 downto 0);
r5: out std_logic_vector(31 downto 0);
r6: out std_logic_vector(31 downto 0);
r7: out std_logic_vector(31 downto 0)
);
end register_file;

architecture bhv of register_file is
type memory is array (0 to 7) of std_logic_vector(31 downto 0);
signal reg: memory;
begin
process(clk,SR1_address,SR2_address,DR_enable, DR_address, data_in)
begin
  if(rst = '1') then
    SR1_out<="00000000000000000000000000000000";
    SR2_out<="00000000000000000000000000000000";
    reg(0)<="00000000000000000000000000000000";
    reg(1)<="00000000000000000000000000000000";
    reg(2)<="00000000000000000000000000000000";
    reg(3)<="00000000000000000000000000000000";
    reg(4)<="00000000000000000000000000000000";
    reg(5)<="00000000000000000000000000000000";
    reg(6)<="00000000000000000000000000000000";
    reg(7)<="00000000000000000000000000000000";
  else
  if(clk'event and clk='1') then
SR1_out <= reg(conv_integer(SR1_address));
SR2_out <= reg(conv_integer(SR2_address));
  if(DR_enable = '1') then
reg(conv_integer(DR_address))<=data_in;
end if;
 end if;
  end if;
end process;

process(clk)
  begin
    r0<= reg(0);
    r1<= reg(1);
    r2<= reg(2);
    r3<= reg(3);
    r4<= reg(4);
    r5<= reg(5);
    r6<= reg(6);
    r7<= reg(7);
  end process;
end bhv;

--LC-2 ALU---------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity LC2_ALU is
port( rst : in std_logic;
A: in std_logic_vector (31 downto 0);
B: in std_logic_vector (31 downto 0);
S: in std_logic; --_vector (1 downto 0);
O: out std_logic_vector (31 downto 0);
EQ: out std_logic);
end LC2_ALU;

architecture bhv of LC2_ALU is
begin
process(A, B, S,rst)
begin
   if(rst ='1') then 
     O<="00000000000000000000000000000000";
     EQ<='0';
   else
case S is
when '0' => O <= A+B;
when '1' => O <= not (A and B);
when others => null;
end case;
if (A=B) then EQ <= '1';
else EQ <= '0';
end if;
end if;
end process;
end bhv;

--controller for the LC-2K?not completed
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
entity FSM is
port(clk: in std_logic;
rst: in std_logic;
OpCode: in std_logic_vector(2 downto 0);
PC_en: out std_logic;
Mem_mux: out std_logic;
Mem_en: out std_logic;
Mem_rw: out std_logic;
IR_en: out std_logic;
Dest_mux: out std_logic;
RData_mux: out std_logic;
Reg_en: out std_logic;
ALU_mux1: out std_logic; --_vector(1 downto 0);
ALU_mux2: out std_logic_vector(1 downto 0);
ALU_op: out std_logic
);
end FSM;


architecture FSM_arch of FSM is
type STATE_TYPE is (FET_0, DEC_1, DEC_2,DEC_3,ADD_4, ADD_5, NAND_6, NAND_7, LW_8, LW_9, LW_10, SW_11, SW_12, BEQ_13, BEQ_14,JALR_15,JALR_16,JALR_17,NOOP_18,HALT_19);
signal cpu_state : STATE_TYPE;
constant ADD : std_logic_vector(2 downto 0) := "000";
constant NAD : std_logic_vector(2 downto 0) := "001";
constant LW : std_logic_vector(2 downto 0) := "010";
constant SW : std_logic_vector(2 downto 0) := "011";
constant BEQ : std_logic_vector(2 downto 0) := "100";
constant JALR : std_logic_vector(2 downto 0) := "101";
constant HALT : std_logic_vector(2 downto 0) := "110";
constant NOOP : std_logic_vector(2 downto 0) := "111";

begin
state_machine : process (rst, clk)
begin
if (rst = '1') then
cpu_state <= FET_0; --reset the controller
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '0';
ALU_mux2 <= "00";
ALU_op <= '0';

elsif (clk'event and clk='1') then
case cpu_state is
--Fetch State---------------------------------------------------------
when FET_0=>
cpu_state <= DEC_1;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '1';
Mem_rw <= '0';
IR_en <= '1';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '0';
ALU_mux2 <= "01";
ALU_op <= '0';

--Decode State---------------------------------------------------------
when DEC_1=>
  cpu_state<= DEC_2;
when DEC_2=>
  cpu_state<=DEC_3;
when DEC_3=>
PC_en <= '1';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '0';
ALU_mux2 <= "01";
ALU_op <= '0';

if (OpCode = ADD ) then
cpu_state <= ADD_4;

elsif (OpCode = NAD ) then
cpu_state <= NAND_6;

elsif (OpCode = LW ) then
cpu_state <= LW_8;

elsif (OpCode = SW ) then
cpu_state <= SW_11;

elsif (OpCode = BEQ ) then
cpu_state <= BEQ_13;

elsif (OpCode = JALR ) then
cpu_state <= JALR_15;

elsif (OpCode = NOOP ) then
cpu_state <= NOOP_18;

elsif (OpCode = HALT ) then
cpu_state <= HALT_19;
end if;

--Add State 4---------------------------------------------------------
when ADD_4=>
cpu_state <= ADD_5;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '1';
ALU_mux2 <= "00";
ALU_op <= '0';

--Add State 5---------------------------------------------------------
when ADD_5=>
cpu_state <= FET_0;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '1';
RData_mux <= '1';
Reg_en <= '1';
ALU_mux1 <= '0';
ALU_mux2 <= "01";
ALU_op <= '0';

--Nand State 6---------------------------------------------------------
when NAND_6=>
cpu_state <= NAND_7;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '1';
ALU_mux2 <= "00";
ALU_op <= '1';

--Nand State 7---------------------------------------------------------
when NAND_7=>
cpu_state <= FET_0;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '1';
RData_mux <= '1';
Reg_en <= '1';
ALU_mux1 <= '0';
ALU_mux2 <= "01";
ALU_op <= '1';

--Load State 8---------------------------------------------------------
when LW_8=>
cpu_state <= LW_9;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '1';
ALU_mux2 <= "11";
ALU_op <= '0';

--Load State 9---------------------------------------------------------
when LW_9=>
cpu_state <= LW_10;
PC_en <= '0';
Mem_mux <= '1';
Mem_en <= '1';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '0';
ALU_mux2 <= "00";
ALU_op <= '0';

--Load State 10---------------------------------------------------------
when LW_10=>
cpu_state <= FET_0;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '1';
ALU_mux1 <= '0';
ALU_mux2 <= "00";
ALU_op <= '0';

--Store State 11---------------------------------------------------------
when SW_11=>
cpu_state <= SW_12;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '1';
ALU_mux2 <= "11";
ALU_op <= '0';

--Store State 12---------------------------------------------------------
when SW_12=>
cpu_state <= FET_0;
PC_en <= '0';
Mem_mux <= '1';
Mem_en <= '1';
Mem_rw <= '1';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '0';
ALU_mux2 <= "00";
ALU_op <= '0';

--branch equal State 13--------------------------------------------------
when BEQ_13=>
cpu_state <= BEQ_14;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '0';
ALU_mux2 <= "11";
ALU_op <= '0';

--branch equal State 14--------------------------------------------------
when BEQ_14=>
cpu_state <= FET_0;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '1';
ALU_mux2 <= "00";
ALU_op <= '0';

--jump register State 15-------------------------------------------------
when JALR_15=>
cpu_state <= JALR_16;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '1';
Reg_en <= '1';
ALU_mux1 <= '0';
ALU_mux2 <= "10";
ALU_op <= '0';

--jump register State 16-------------------------------------------------
when JALR_16=>
cpu_state <= JALR_17;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '1';
ALU_mux2 <= "10";
ALU_op <= '0';
--jump register State 17-------------------------------------------------
when JALR_17=>
cpu_state <= FET_0;
PC_en <= '1';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '1';
ALU_mux2 <= "10";
ALU_op <= '0';

--no operation 18--------------------------------------------------------
when NOOP_18=>
cpu_state <= FET_0;

--halt State 19----------------------------------------------------------
when HALT_19=>
cpu_state <= HALT_19;
PC_en <= '0';
Mem_mux <= '0';
Mem_en <= '0';
Mem_rw <= '0';
IR_en <= '0';
Dest_mux <= '0';
RData_mux <= '0';
Reg_en <= '0';
ALU_mux1 <= '0';
ALU_mux2 <= "00";
ALU_op <= '0';

---------------------------------------------------------------------
end case;
end if;
end process state_machine;
end FSM_arch;

--Datapath and Controller combined structurally---------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity LC2_all is
port(rst: in STD_LOGIC;
clk: in STD_LOGIC);
end LC2_all;

architecture str of LC2_all is
  
component LC2_ALU
port( rst: in std_logic;
A: in std_logic_vector (31 downto 0);
B: in std_logic_vector (31 downto 0);
S: in std_logic; --_vector (1 downto 0);
O: out std_logic_vector (31 downto 0);
EQ: out std_logic);
end component;

component branch
 port(rst :in std_logic;
    beq :in std_logic;
    opcode :in std_logic_vector(2 downto 0);
    pccontrol :in std_logic;
    pcen:out std_logic);
end component;

component muxr
port(rst: in std_logic;
c : in std_logic_vector(2 downto 0);
d : in std_logic_vector(2 downto 0);
s : in std_logic;
muxoutput : out std_logic_vector(2 downto 0));
end component;

component mux2
port(rst: std_logic;
c : in std_logic_vector(31 downto 0);
d : in std_logic_vector(31 downto 0);
s : in std_logic;
muxoutput : out std_logic_vector(31 downto 0));
end component;

component mux4
port(rst : std_logic;
c : in std_logic_vector(31 downto 0);
d : in std_logic_vector(31 downto 0);
e : in std_logic_vector(31 downto 0);
f : in std_logic_vector(31 downto 0);
s : in std_logic_vector(1 downto 0);
muxoutput : out std_logic_vector(31 downto 0));
end component;

component reg
port(rst :std_logic;
clk : in std_logic;
enable : in std_logic;
data : in std_logic_vector (31 downto 0);
O : out std_logic_vector (31 downto 0));
end component;

component register_file
port(rst :std_logic;
clk : in std_logic;
DR_enable : in std_logic;
DR_address : in std_logic_vector (2 downto 0);
SR1_address: in std_logic_vector(2 downto 0);
SR2_address: in std_logic_vector(2 downto 0);
data_in: in std_logic_vector (31 downto 0);
SR1_out: out std_logic_vector (31 downto 0);
SR2_out: out std_logic_vector (31 downto 0);
r0: out std_logic_vector(31 downto 0);
r1: out std_logic_vector(31 downto 0);
r2: out std_logic_vector(31 downto 0);
r3: out std_logic_vector(31 downto 0);
r4: out std_logic_vector(31 downto 0);
r5: out std_logic_vector(31 downto 0);
r6: out std_logic_vector(31 downto 0);
r7: out std_logic_vector(31 downto 0)
);
end component;

component sext
port(rst :std_logic;
A : in std_logic_vector (15 downto 0);
O : out std_logic_vector (31 downto 0));
end component;

component ram_module
port(rst : in std_logic;
clk : in std_logic;
enable : in std_logic;
R_W : in std_logic;
addr : in std_logic_vector (31 downto 0);
data_in : in std_logic_vector (31 downto 0);
data_out : out std_logic_vector (31 downto 0));
end component;

component FSM
port(clk: in std_logic;
rst: in std_logic;
OpCode: in std_logic_vector(2 downto 0);
PC_en: out std_logic;
Mem_mux: out std_logic;
Mem_en: out std_logic;
Mem_rw: out std_logic;
IR_en: out std_logic;
Dest_mux: out std_logic;
RData_mux: out std_logic;
Reg_en: out std_logic;
ALU_mux1: out std_logic; --_vector(1 downto 0);
ALU_mux2: out std_logic_vector(1 downto 0);
ALU_op: out std_logic);
end component;

signal PCout : std_logic_vector(31 downto 0);
signal ALUresult : std_logic_vector(31 downto 0);
signal PCen : std_logic;
signal PCBRANCHen: std_logic ;
signal ADDRout : std_logic_vector(31 downto 0);
signal ADDRmux : std_logic;
signal RAMout : std_logic_vector(31 downto 0);
signal MEMen : std_logic;
signal RW : std_logic;
signal IRout : std_logic_vector(31 downto 0);
signal IRen : std_logic;
signal REGW : std_logic_vector(2 downto 0);
signal REGdata : std_logic_vector(31 downto 0);
signal DESTmux : std_logic;
signal REGmux2 : std_logic;
signal REGen : std_logic;
signal REGout1 : std_logic_vector(31 downto 0);
signal REGout2 : std_logic_vector(31 downto 0);
signal SEXTout : std_logic_vector(31 downto 0);
signal ALU1 : std_logic_vector(31 downto 0);
signal ALU2 : std_logic_vector(31 downto 0);
signal ALUmux1 : std_logic;
signal ALUmux2 : std_logic_vector(1 downto 0);
signal ALUout : std_logic_vector(31 downto 0);
signal ALUsel : std_logic;
signal ALUeql :std_logic;
signal ground : std_logic;
signal ground32 : std_logic_vector(31 downto 0);
signal Vcc : std_logic;
signal r0:std_logic_vector(31 downto 0):= "00000000000000000000000000000000";
signal r1:std_logic_vector(31 downto 0):= "00000000000000000000000000000000";
signal r2:std_logic_vector(31 downto 0):= "00000000000000000000000000000000";
signal r3:std_logic_vector(31 downto 0):= "00000000000000000000000000000000";
signal r4:std_logic_vector(31 downto 0):= "00000000000000000000000000000000";
signal r5:std_logic_vector(31 downto 0):= "00000000000000000000000000000000";
signal r6:std_logic_vector(31 downto 0):= "00000000000000000000000000000000";
signal r7:std_logic_vector(31 downto 0):= "00000000000000000000000000000000";


begin
ground <= '0';
ground32 <= "00000000000000000000000000000000";
Vcc <= '1';

U_PC : reg port map (rst,clk, PCBRANCHen , ALUresult,PCout);
U_ADDR_mux : mux2 port map (rst,PCout, ALUresult, ADDRmux, ADDRout);
U_ram : ram_module port map (rst,clk, MEMen, RW, ADDRout, REGout2, RAMout);
U_IR_reg : reg port map (rst,clk, IRen, RAMout, IRout);
U_FSM : FSM port map (clk, rst, IRout(24 downto 22), PCen,ADDRmux, MEMen,RW, IRen,DESTmux,REGmux2,REGen, ALUmux1, ALUmux2, ALUsel);
U_REG_mux1 : muxr port map (rst,IRout(18 downto 16), IRout(2 downto 0), DESTmux, REGW(2 downto 0));
U_REG_mux2 : mux2 port map (rst,RAMout, ALUresult, REGmux2, REGdata);
U_REG_bank : register_file port map (rst,clk, REGen, REGW, IRout(21 downto 19), IRout(18 downto 16), REGdata, REGout1, REGout2,r0,r1,
r2,r3,r4,r5,r6,r7);
U_sext : sext port map (rst,IRout(15 downto 0), SEXTout);
U_ALU_mux1 : mux2 port map (rst,PCout, REGout1, ALUmux1, ALU1);
U_ALU_mux2 : mux4 port map (rst,REGout2, conv_std_logic_vector(1,32),conv_std_logic_vector(0,32),SEXTout, ALUmux2, ALU2);
U_ALU : LC2_ALU port map (rst,ALU1, ALU2,ALUsel,ALUout, ALUeql);
U_PC_BRANCH_EN: branch port map(rst,ALUeql,IRout(24 downto 22),PCen,PCBRANCHen);
U_ALU_reg : reg port map (rst,clk, Vcc, ALUout, ALUresult); 
end str;


--Test bench--------------------------------------------------

library ieee;
use ieee.std_logic_arith.all;
use ieee.STD_LOGIC_UNSIGNED.all;
use ieee.std_logic_1164.all;

-- Add your library and packages declaration here ...
entity lc2_all_tb is
end lc2_all_tb;

architecture TB_ARCHITECTURE of lc2_all_tb is
-- Component declaration of the tested unit
component LC2_all
port(
rst : in std_logic;
clk : in std_logic );
end component;

-- Stimulus signals - signals mapped to the input and inout ports of tested
signal rst : std_logic:='1';
signal clk : std_logic;
-- Observed signals - signals mapped to the output ports of tested entity
begin
-- Unit Under Test port map 
process
begin
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
end process; 

process
begin
rst <= '0' after 1 ns;
wait;
end process;

UUT : LC2_all port map(rst,clk);
end TB_ARCHITECTURE;

configuration TESTBENCH_FOR_LC2_all of lc2_all_tb is
for TB_ARCHITECTURE
for UUT : LC2_all
use entity work.LC2_all(str);
end for;
end for;
end TESTBENCH_FOR_LC2_all;

